LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

--Component that maps acceleration to angle

ENTITY angle_converter IS
    PORT (
        in_val :  IN INTEGER;    --acceleration in either the X or the Y axis. In range 0-128
        z_MSB  :  IN STD_LOGIC;  --MSB av accelerationen i Z-öed
        angle  :  OUT INTEGER    --Outputs the angle
    );
END angle_converter;



ARCHITECTURE Behavioral OF angle_converter IS

    BEGIN
        PROCESS(in_val, z_MSB)
        --Maps the interval 0-129 to 0-90 degrees
        --To find what values that maps to what angle we used this formila:
        --       y = round_off(x * 90/129)
        --Where x is the in_val and y is the corresponding angle
            BEGIN
                IF z_MSB = '0' THEN       
                    CASE in_val IS
                        WHEN 0 => angle <= 0;
                        WHEN 1 => angle <= 1;
                        WHEN 2 => angle <= 1;
                        WHEN 3 => angle <= 2;
                        WHEN 4 => angle <= 3;
                        WHEN 5 => angle <= 3;
                        WHEN 6 => angle <= 4;
                        WHEN 7 => angle <= 5;
                        WHEN 8 => angle <= 6;
                        WHEN 9 => angle <= 6;
                        WHEN 10 => angle <= 7;
                        WHEN 11 => angle <= 8;
                        WHEN 12 => angle <= 8;
                        WHEN 13 => angle <= 9;
                        WHEN 14 => angle <= 10;
                        WHEN 15 => angle <= 10;
                        WHEN 16 => angle <= 11;
                        WHEN 17 => angle <= 12;
                        WHEN 18 => angle <= 12;
                        WHEN 19 => angle <= 13;
                        WHEN 20 => angle <= 14;
                        WHEN 21 => angle <= 15;
                        WHEN 22 => angle <= 15;
                        WHEN 23 => angle <= 16;
                        WHEN 24 => angle <= 17;
                        WHEN 25 => angle <= 17;
                        WHEN 26 => angle <= 18;
                        WHEN 27 => angle <= 19;
                        WHEN 28 => angle <= 19;
                        WHEN 29 => angle <= 20;
                        WHEN 30 => angle <= 21;
                        WHEN 31 => angle <= 21;
                        WHEN 32 => angle <= 22;
                        WHEN 33 => angle <= 23;
                        WHEN 34 => angle <= 24;
                        WHEN 35 => angle <= 24;
                        WHEN 36 => angle <= 25;
                        WHEN 37 => angle <= 26;
                        WHEN 38 => angle <= 26;
                        WHEN 39 => angle <= 27;
                        WHEN 40 => angle <= 28;
                        WHEN 41 => angle <= 28;
                        WHEN 42 => angle <= 29;
                        WHEN 43 => angle <= 30;
                        WHEN 44 => angle <= 30;
                        WHEN 45 => angle <= 31;
                        WHEN 46 => angle <= 32;
                        WHEN 47 => angle <= 33;
                        WHEN 48 => angle <= 33;
                        WHEN 49 => angle <= 34;
                        WHEN 50 => angle <= 35;
                        WHEN 51 => angle <= 35;
                        WHEN 52 => angle <= 36;
                        WHEN 53 => angle <= 37;
                        WHEN 54 => angle <= 37;
                        WHEN 55 => angle <= 38;
                        WHEN 56 => angle <= 39;
                        WHEN 57 => angle <= 39;
                        WHEN 58 => angle <= 40;
                        WHEN 59 => angle <= 41;
                        WHEN 60 => angle <= 42;
                        WHEN 61 => angle <= 42;
                        WHEN 62 => angle <= 43;
                        WHEN 63 => angle <= 44;
                        WHEN 64 => angle <= 44;
                        WHEN 65 => angle <= 45;
                        WHEN 66 => angle <= 46;
                        WHEN 67 => angle <= 46;
                        WHEN 68 => angle <= 47;
                        WHEN 69 => angle <= 48;
                        WHEN 70 => angle <= 48;
                        WHEN 71 => angle <= 49;
                        WHEN 72 => angle <= 50;
                        WHEN 73 => angle <= 51;
                        WHEN 74 => angle <= 51;
                        WHEN 75 => angle <= 52;
                        WHEN 76 => angle <= 53;
                        WHEN 77 => angle <= 53;
                        WHEN 78 => angle <= 54;
                        WHEN 79 => angle <= 55;
                        WHEN 80 => angle <= 55;
                        WHEN 81 => angle <= 56;
                        WHEN 82 => angle <= 57;
                        WHEN 83 => angle <= 57;
                        WHEN 84 => angle <= 58;
                        WHEN 85 => angle <= 59;
                        WHEN 86 => angle <= 60;
                        WHEN 87 => angle <= 60;
                        WHEN 88 => angle <= 61;
                        WHEN 89 => angle <= 62;
                        WHEN 90 => angle <= 62;
                        WHEN 91 => angle <= 63;
                        WHEN 92 => angle <= 64;
                        WHEN 93 => angle <= 64;
                        WHEN 94 => angle <= 65;
                        WHEN 95 => angle <= 66;
                        WHEN 96 => angle <= 66;
                        WHEN 97 => angle <= 67;
                        WHEN 98 => angle <= 68;
                        WHEN 99 => angle <= 69;
                        WHEN 100 => angle <= 69;
                        WHEN 101 => angle <= 70;
                        WHEN 102 => angle <= 71;
                        WHEN 103 => angle <= 71;
                        WHEN 104 => angle <= 72;
                        WHEN 105 => angle <= 73;
                        WHEN 106 => angle <= 73;
                        WHEN 107 => angle <= 74;
                        WHEN 108 => angle <= 75;
                        WHEN 109 => angle <= 75;
                        WHEN 110 => angle <= 76;
                        WHEN 111 => angle <= 77;
                        WHEN 112 => angle <= 78;
                        WHEN 113 => angle <= 78;
                        WHEN 114 => angle <= 79;
                        WHEN 115 => angle <= 80;
                        WHEN 116 => angle <= 80;
                        WHEN 117 => angle <= 81;
                        WHEN 118 => angle <= 82;
                        WHEN 119 => angle <= 82;
                        WHEN 120 => angle <= 83;
                        WHEN 121 => angle <= 84;
                        WHEN 122 => angle <= 84;
                        WHEN 123 => angle <= 85;
                        WHEN 124 => angle <= 86;
                        WHEN 125 => angle <= 87;
                        WHEN 126 => angle <= 87;
                        WHEN 127 => angle <= 88;
                        WHEN 128 => angle <= 89;
                        WHEN 129 => angle <= 90;
                        WHEN OTHERS => angle <= 90;
                     END CASE;
                ELSE
                --Angles when MSB(Z) = '1'
                --This means that the spirit level is leaning >90 degrees
                    CASE in_val IS
                        WHEN 0 => angle <= 180-0;
                        WHEN 1 => angle <= 180-1;
                        WHEN 2 => angle <= 180-1;
                        WHEN 3 => angle <= 180-2;
                        WHEN 4 => angle <= 180-3;
                        WHEN 5 => angle <= 180-3;
                        WHEN 6 => angle <= 180-4;
                        WHEN 7 => angle <= 180-5;
                        WHEN 8 => angle <= 180-6;
                        WHEN 9 => angle <= 180-6;
                        WHEN 10 => angle <= 180-7;
                        WHEN 11 => angle <= 180-8;
                        WHEN 12 => angle <= 180-8;
                        WHEN 13 => angle <= 180-9;
                        WHEN 14 => angle <= 180-10;
                        WHEN 15 => angle <= 180-10;
                        WHEN 16 => angle <= 180-11;
                        WHEN 17 => angle <= 180-12;
                        WHEN 18 => angle <= 180-12;
                        WHEN 19 => angle <= 180-13;
                        WHEN 20 => angle <= 180-14;
                        WHEN 21 => angle <= 180-15;
                        WHEN 22 => angle <= 180-15;
                        WHEN 23 => angle <= 180-16;
                        WHEN 24 => angle <= 180-17;
                        WHEN 25 => angle <= 180-17;
                        WHEN 26 => angle <= 180-18;
                        WHEN 27 => angle <= 180-19;
                        WHEN 28 => angle <= 180-19;
                        WHEN 29 => angle <= 180-20;
                        WHEN 30 => angle <= 180-21;
                        WHEN 31 => angle <= 180-21;
                        WHEN 32 => angle <= 180-22;
                        WHEN 33 => angle <= 180-23;
                        WHEN 34 => angle <= 180-24;
                        WHEN 35 => angle <= 180-24;
                        WHEN 36 => angle <= 180-25;
                        WHEN 37 => angle <= 180-26;
                        WHEN 38 => angle <= 180-26;
                        WHEN 39 => angle <= 180-27;
                        WHEN 40 => angle <= 180-28;
                        WHEN 41 => angle <= 180-28;
                        WHEN 42 => angle <= 180-29;
                        WHEN 43 => angle <= 180-30;
                        WHEN 44 => angle <= 180-30;
                        WHEN 45 => angle <= 180-31;
                        WHEN 46 => angle <= 180-32;
                        WHEN 47 => angle <= 180-33;
                        WHEN 48 => angle <= 180-33;
                        WHEN 49 => angle <= 180-34;
                        WHEN 50 => angle <= 180-35;
                        WHEN 51 => angle <= 180-35;
                        WHEN 52 => angle <= 180-36;
                        WHEN 53 => angle <= 180-37;
                        WHEN 54 => angle <= 180-37;
                        WHEN 55 => angle <= 180-38;
                        WHEN 56 => angle <= 180-39;
                        WHEN 57 => angle <= 180-39;
                        WHEN 58 => angle <= 180-40;
                        WHEN 59 => angle <= 180-41;
                        WHEN 60 => angle <= 180-42;
                        WHEN 61 => angle <= 180-42;
                        WHEN 62 => angle <= 180-43;
                        WHEN 63 => angle <= 180-44;
                        WHEN 64 => angle <= 180-44;
                        WHEN 65 => angle <= 180-45;
                        WHEN 66 => angle <= 180-46;
                        WHEN 67 => angle <= 180-46;
                        WHEN 68 => angle <= 180-47;
                        WHEN 69 => angle <= 180-48;
                        WHEN 70 => angle <= 180-48;
                        WHEN 71 => angle <= 180-49;
                        WHEN 72 => angle <= 180-50;
                        WHEN 73 => angle <= 180-51;
                        WHEN 74 => angle <= 180-51;
                        WHEN 75 => angle <= 180-52;
                        WHEN 76 => angle <= 180-53;
                        WHEN 77 => angle <= 180-53;
                        WHEN 78 => angle <= 180-54;
                        WHEN 79 => angle <= 180-55;
                        WHEN 80 => angle <= 180-55;
                        WHEN 81 => angle <= 180-56;
                        WHEN 82 => angle <= 180-57;
                        WHEN 83 => angle <= 180-57;
                        WHEN 84 => angle <= 180-58;
                        WHEN 85 => angle <= 180-59;
                        WHEN 86 => angle <= 180-60;
                        WHEN 87 => angle <= 180-60;
                        WHEN 88 => angle <= 180-61;
                        WHEN 89 => angle <= 180-62;
                        WHEN 90 => angle <= 180-62;
                        WHEN 91 => angle <= 180-63;
                        WHEN 92 => angle <= 180-64;
                        WHEN 93 => angle <= 180-64;
                        WHEN 94 => angle <= 180-65;
                        WHEN 95 => angle <= 180-66;
                        WHEN 96 => angle <= 180-66;
                        WHEN 97 => angle <= 180-67;
                        WHEN 98 => angle <= 180-68;
                        WHEN 99 => angle <= 180-69;
                        WHEN 100 => angle <= 180-69;
                        WHEN 101 => angle <= 180-70;
                        WHEN 102 => angle <= 180-71;
                        WHEN 103 => angle <= 180-71;
                        WHEN 104 => angle <= 180-72;
                        WHEN 105 => angle <= 180-73;
                        WHEN 106 => angle <= 180-73;
                        WHEN 107 => angle <= 180-74;
                        WHEN 108 => angle <= 180-75;
                        WHEN 109 => angle <= 180-75;
                        WHEN 110 => angle <= 180-76;
                        WHEN 111 => angle <= 180-77;
                        WHEN 112 => angle <= 180-78;
                        WHEN 113 => angle <= 180-78;
                        WHEN 114 => angle <= 180-79;
                        WHEN 115 => angle <= 180-80;
                        WHEN 116 => angle <= 180-80;
                        WHEN 117 => angle <= 180-81;
                        WHEN 118 => angle <= 180-82;
                        WHEN 119 => angle <= 180-82;
                        WHEN 120 => angle <= 180-83;
                        WHEN 121 => angle <= 180-84;
                        WHEN 122 => angle <= 180-84;
                        WHEN 123 => angle <= 180-85;
                        WHEN 124 => angle <= 180-86;
                        WHEN 125 => angle <= 180-87;
                        WHEN 126 => angle <= 180-87;
                        WHEN 127 => angle <= 180-88;
                        WHEN 128 => angle <= 180-89;
                        WHEN 129 => angle <= 180-89;
                        WHEN OTHERS => angle <= 180-90;
                     END CASE;
            END IF;
    END PROCESS; 
END Behavioral;
